module N_bit_Adder_Subtractor (
    ports
);
    
endmodule






