module and (
    out, in1, in2
) (
    input in1, in2;
    output out;
);
    
endmodule